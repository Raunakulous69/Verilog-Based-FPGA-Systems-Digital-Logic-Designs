module hex7seg
(
   input [3:0] N,
   
   output [6:0] Seg
);
  
  assign Seg[0] = (~N[3]&~N[2]&~N[1]&N[0])|(~N[3]&N[2]&~N[1]&~N[0])|(N[3]&~N[2]&N[1]&N[0])|(N[3]&N[2]&~N[1]&N[0]);
  assign Seg[1] = (~N[3]&N[2]&~N[1]&N[0])|(~N[3]&N[2]&N[1]&~N[0])|(N[3]&~N[2]&N[1]&N[0])|(N[3]&N[2]&~N[1]&~N[0])|(N[3]&N[2]&N[1]&~N[0])|(N[3]&N[2]&N[1]&N[0]);
  assign Seg[2] = (~N[3]&~N[2]&N[1]&~N[0])|(N[3]&N[2]&~N[1]&~N[0])|(N[3]&N[2]&N[1]&~N[0])|(N[3]&N[2]&N[1]&N[0]);
  assign Seg[3] = (~N[3]&~N[2]&~N[1]&N[0])|(~N[3]&N[2]&~N[1]&~N[0])|(~N[3]&N[2]&N[1]&N[0])|(N[3]&~N[2]&~N[1]&N[0])|(N[3]&~N[2]&N[1]&~N[0])|(N[3]&N[2]&N[1]&N[0]);
  assign Seg[4] = (~N[3]&~N[2]&~N[1]&N[0])|(~N[3]&~N[2]&N[1]&N[0])|(~N[3]&N[2]&~N[1]&~N[0])|(~N[3]&N[2]&~N[1]&N[0])|(~N[3]&N[2]&N[1]&N[0])|(N[3]&~N[2]&~N[1]&N[0]);
  assign Seg[5] = (~N[3]&~N[2]&~N[1]&N[0])|(~N[3]&~N[2]&N[1]&~N[0])|(~N[3]&~N[2]&N[1]&N[0])|(~N[3]&N[2]&N[1]&N[0])|(N[3]&N[2]&~N[1]&N[0]);
  assign Seg[6] = (~N[3]&~N[2]&~N[1]&~N[0])|(~N[3]&~N[2]&~N[1]&N[0])|(~N[3]&N[2]&N[1]&N[0])|(N[3]&N[2]&~N[1]&~N[0]);
 
endmodule

